class fifo_sbd extends uvm_scoreboard;

`uvm_component_utils(fifo_sbd)
function new(string name,uvm_component parent);
	super.new(name,parent);
endfunction
endclass

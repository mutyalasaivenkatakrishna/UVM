
typedef uvm_sequencer#(fifo_tx) fifo_sqr;

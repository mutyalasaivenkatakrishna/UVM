`define DEPTH 10
`define WIDTH 10
`define AD_W $clog2(DEPTH)



